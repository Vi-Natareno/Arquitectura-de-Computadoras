//Definicion del modulo y sus i/p
module _and (input A, input B, output C); //puede comenzar solo con guion bajo, mayus o minus
//2. declara señales/ elementos internos


//3. Comportamiento del modulo 
//(asignaciones, instancias, conexiones)
//
assign C = A&B;
 
 
 endmodule